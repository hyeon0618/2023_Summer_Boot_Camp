library verilog;
use verilog.vl_types.all;
entity tb_ring is
end tb_ring;
