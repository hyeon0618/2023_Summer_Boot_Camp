module alu (
    input clk,
    input n_rst,
    input [3:0] dtype,
    input [4:0] operator,
    input parser_done,
    input [31:0] src1, src2,
    output alu_done,
    output calc_res
);
    
endmodule