library verilog;
use verilog.vl_types.all;
entity tb_d_ff is
end tb_d_ff;
