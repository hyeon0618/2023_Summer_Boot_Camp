module decoder (
    input clk,
    input n_rst,
    input [7:0] data,
    input dout_valid,
    output [3:0] data_type,
    output [4:0] operator,
    output parser_done,
    output [31:0] src1, src2
);


    
endmodule