library verilog;
use verilog.vl_types.all;
entity test is
    port(
        a               : in     vl_logic;
        \out\           : out    vl_logic
    );
end test;
