module encoder (
    input clk,
    input n_rst,
    input alu_done,
    input [31:0] result,
    input uin_ready,
    output [7:0] uart_out,
    output uout_valid
);
    
endmodule